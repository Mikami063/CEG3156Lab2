library verilog;
use verilog.vl_types.all;
entity RegsiterFIleTest_vlg_vec_tst is
end RegsiterFIleTest_vlg_vec_tst;
